library verilog;
use verilog.vl_types.all;
entity tb_parking_controller is
end tb_parking_controller;
